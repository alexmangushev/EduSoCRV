library verilog;
use verilog.vl_types.all;
entity gpio_tb is
end gpio_tb;
