import core_pkg::*;
module load_store_unit
(
   input  logic                  clk,
	input  logic                  mem_op,
	input  logic [ADDR_WIDTH-1:0] rd_addr
);
endmodule