package core_pkg;
  parameter    INSTR_WIDTH    = 32; // Instruction width             
  parameter    DATA_WIDTH     = 32; // Data width
  parameter    REG_WIDTH      = 32; // General purpose register width
  parameter    ADDR_WIDTH     = 32; // Address width 
endpackage